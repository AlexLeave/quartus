module _74ls148(I, Y, )



endmodule