library verilog;
use verilog.vl_types.all;
entity keshe_vlg_vec_tst is
end keshe_vlg_vec_tst;
