module des_signal(arr, des_floor)
input arr;
output des_floor;




endmodule