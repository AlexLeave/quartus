module out_3(clk, p);
inout p;
input clk;

reg p;
always@ (negedge clk)
;

endmodule